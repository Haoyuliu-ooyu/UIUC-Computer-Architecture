module keypad(valid, number, a, b, c, d, e, f, g);
   output 	valid;
   output [3:0] number;
   input 	a, b, c, d, e, f, g;
   wire w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, wb0, wb1, wb2, wb3;
   and a0(w0, b, g);
   and a1(w1, a, d);
   and a2(w2, b, d);
   and a3(w3, c, d);
   and a4(w4, a, e);
   and a5(w5, b, e);
   and a6(w6, c, e);
   and a7(w7, a, f);
   and a8(w8, b, f);
   and a9(w9, c, f);
   or o1(valid, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9);
   or o2(wb0, w1, w3, w5, w7, w9);
   or o3(wb1, w2, w3, w6, w7);
   or o4(wb2, w4, w5, w6, w7);
   or o5(wb3, w8, w9);
   assign number[0] = wb0;
   assign number[1] = wb1;
   assign number[2] = wb2;
   assign number[3] = wb3;
endmodule // keypad
